package prog1;

	module mkprog1(Empty);
	
		rule rl_1;
			$display("Hello world");
			$finish(0);
		endrule
	endmodule
endpackage
